library verilog;
use verilog.vl_types.all;
entity testbench_mips is
end testbench_mips;
